module Sort4( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  input  [15:0] io_in0, // @[:@6.4]
  input  [15:0] io_in1, // @[:@6.4]
  input  [15:0] io_in2, // @[:@6.4]
  input  [15:0] io_in3, // @[:@6.4]
  output [15:0] io_out0, // @[:@6.4]
  output [15:0] io_out1, // @[:@6.4]
  output [15:0] io_out2, // @[:@6.4]
  output [15:0] io_out3 // @[:@6.4]
);
  wire  _T_25; // @[Sort4.scala 21:15:@12.4]
  wire [15:0] row10; // @[Sort4.scala 21:25:@13.4]
  wire [15:0] row11; // @[Sort4.scala 21:25:@13.4]
  wire  _T_26; // @[Sort4.scala 29:15:@21.4]
  wire [15:0] row12; // @[Sort4.scala 29:25:@22.4]
  wire [15:0] row13; // @[Sort4.scala 29:25:@22.4]
  wire  _T_29; // @[Sort4.scala 40:14:@32.4]
  wire [15:0] row21; // @[Sort4.scala 40:23:@33.4]
  wire [15:0] row22; // @[Sort4.scala 40:23:@33.4]
  wire  _T_32; // @[Sort4.scala 50:14:@43.4]
  wire [15:0] row20; // @[Sort4.scala 50:23:@44.4]
  wire [15:0] row23; // @[Sort4.scala 50:23:@44.4]
  wire  _T_33; // @[Sort4.scala 58:14:@52.4]
  wire  _T_34; // @[Sort4.scala 66:14:@61.4]
  assign _T_25 = io_in0 < io_in1; // @[Sort4.scala 21:15:@12.4]
  assign row10 = _T_25 ? io_in0 : io_in1; // @[Sort4.scala 21:25:@13.4]
  assign row11 = _T_25 ? io_in1 : io_in0; // @[Sort4.scala 21:25:@13.4]
  assign _T_26 = io_in2 < io_in3; // @[Sort4.scala 29:15:@21.4]
  assign row12 = _T_26 ? io_in2 : io_in3; // @[Sort4.scala 29:25:@22.4]
  assign row13 = _T_26 ? io_in3 : io_in2; // @[Sort4.scala 29:25:@22.4]
  assign _T_29 = row11 < row12; // @[Sort4.scala 40:14:@32.4]
  assign row21 = _T_29 ? row11 : row12; // @[Sort4.scala 40:23:@33.4]
  assign row22 = _T_29 ? row12 : row11; // @[Sort4.scala 40:23:@33.4]
  assign _T_32 = row10 < row13; // @[Sort4.scala 50:14:@43.4]
  assign row20 = _T_32 ? row10 : row13; // @[Sort4.scala 50:23:@44.4]
  assign row23 = _T_32 ? row13 : row10; // @[Sort4.scala 50:23:@44.4]
  assign _T_33 = row20 < row21; // @[Sort4.scala 58:14:@52.4]
  assign _T_34 = row22 < row23; // @[Sort4.scala 66:14:@61.4]
  assign io_out0 = _T_33 ? row20 : row21; // @[Sort4.scala 59:13:@54.6 Sort4.scala 62:13:@58.6]
  assign io_out1 = _T_33 ? row21 : row20; // @[Sort4.scala 60:13:@55.6 Sort4.scala 63:13:@59.6]
  assign io_out2 = _T_34 ? row22 : row23; // @[Sort4.scala 67:13:@63.6 Sort4.scala 70:13:@67.6]
  assign io_out3 = _T_34 ? row23 : row22; // @[Sort4.scala 68:13:@64.6 Sort4.scala 71:13:@68.6]
endmodule
