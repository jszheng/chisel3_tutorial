module MaxN( // @[:@3.2]
  input        clock, // @[:@4.4]
  input        reset, // @[:@5.4]
  input  [7:0] io_ins_0, // @[:@6.4]
  input  [7:0] io_ins_1, // @[:@6.4]
  input  [7:0] io_ins_2, // @[:@6.4]
  input  [7:0] io_ins_3, // @[:@6.4]
  input  [7:0] io_ins_4, // @[:@6.4]
  input  [7:0] io_ins_5, // @[:@6.4]
  input  [7:0] io_ins_6, // @[:@6.4]
  input  [7:0] io_ins_7, // @[:@6.4]
  input  [7:0] io_ins_8, // @[:@6.4]
  input  [7:0] io_ins_9, // @[:@6.4]
  output [7:0] io_out // @[:@6.4]
);
  wire  _T_37; // @[MaxN.scala 10:46:@8.4]
  wire [7:0] _T_38; // @[MaxN.scala 10:43:@9.4]
  wire  _T_39; // @[MaxN.scala 10:46:@10.4]
  wire [7:0] _T_40; // @[MaxN.scala 10:43:@11.4]
  wire  _T_41; // @[MaxN.scala 10:46:@12.4]
  wire [7:0] _T_42; // @[MaxN.scala 10:43:@13.4]
  wire  _T_43; // @[MaxN.scala 10:46:@14.4]
  wire [7:0] _T_44; // @[MaxN.scala 10:43:@15.4]
  wire  _T_45; // @[MaxN.scala 10:46:@16.4]
  wire [7:0] _T_46; // @[MaxN.scala 10:43:@17.4]
  wire  _T_47; // @[MaxN.scala 10:46:@18.4]
  wire [7:0] _T_48; // @[MaxN.scala 10:43:@19.4]
  wire  _T_49; // @[MaxN.scala 10:46:@20.4]
  wire [7:0] _T_50; // @[MaxN.scala 10:43:@21.4]
  wire  _T_51; // @[MaxN.scala 10:46:@22.4]
  wire [7:0] _T_52; // @[MaxN.scala 10:43:@23.4]
  wire  _T_53; // @[MaxN.scala 10:46:@24.4]
  assign _T_37 = io_ins_0 > io_ins_1; // @[MaxN.scala 10:46:@8.4]
  assign _T_38 = _T_37 ? io_ins_0 : io_ins_1; // @[MaxN.scala 10:43:@9.4]
  assign _T_39 = _T_38 > io_ins_2; // @[MaxN.scala 10:46:@10.4]
  assign _T_40 = _T_39 ? _T_38 : io_ins_2; // @[MaxN.scala 10:43:@11.4]
  assign _T_41 = _T_40 > io_ins_3; // @[MaxN.scala 10:46:@12.4]
  assign _T_42 = _T_41 ? _T_40 : io_ins_3; // @[MaxN.scala 10:43:@13.4]
  assign _T_43 = _T_42 > io_ins_4; // @[MaxN.scala 10:46:@14.4]
  assign _T_44 = _T_43 ? _T_42 : io_ins_4; // @[MaxN.scala 10:43:@15.4]
  assign _T_45 = _T_44 > io_ins_5; // @[MaxN.scala 10:46:@16.4]
  assign _T_46 = _T_45 ? _T_44 : io_ins_5; // @[MaxN.scala 10:43:@17.4]
  assign _T_47 = _T_46 > io_ins_6; // @[MaxN.scala 10:46:@18.4]
  assign _T_48 = _T_47 ? _T_46 : io_ins_6; // @[MaxN.scala 10:43:@19.4]
  assign _T_49 = _T_48 > io_ins_7; // @[MaxN.scala 10:46:@20.4]
  assign _T_50 = _T_49 ? _T_48 : io_ins_7; // @[MaxN.scala 10:43:@21.4]
  assign _T_51 = _T_50 > io_ins_8; // @[MaxN.scala 10:46:@22.4]
  assign _T_52 = _T_51 ? _T_50 : io_ins_8; // @[MaxN.scala 10:43:@23.4]
  assign _T_53 = _T_52 > io_ins_9; // @[MaxN.scala 10:46:@24.4]
  assign io_out = _T_53 ? _T_52 : io_ins_9; // @[MaxN.scala 16:10:@26.4]
endmodule
