module MyOperators( // @[:@3.2]
  input        clock, // @[:@4.4]
  input        reset, // @[:@5.4]
  input  [3:0] io_in, // @[:@6.4]
  output [3:0] io_out_add, // @[:@6.4]
  output [3:0] io_out_sub, // @[:@6.4]
  output [3:0] io_out_mul // @[:@6.4]
);
  wire [2:0] _T_19; // @[MyOperators.scala 12:21:@11.4]
  wire [2:0] _T_20; // @[MyOperators.scala 12:21:@12.4]
  wire [1:0] _T_21; // @[MyOperators.scala 12:21:@13.4]
  wire [4:0] _T_24; // @[MyOperators.scala 13:21:@15.4]
  assign _T_19 = 2'h2 - 2'h1; // @[MyOperators.scala 12:21:@11.4]
  assign _T_20 = $unsigned(_T_19); // @[MyOperators.scala 12:21:@12.4]
  assign _T_21 = _T_20[1:0]; // @[MyOperators.scala 12:21:@13.4]
  assign _T_24 = 3'h4 * 3'h2; // @[MyOperators.scala 13:21:@15.4]
  assign io_out_add = 4'h5; // @[MyOperators.scala 11:14:@10.4]
  assign io_out_sub = {{2'd0}, _T_21}; // @[MyOperators.scala 12:14:@14.4]
  assign io_out_mul = _T_24[3:0]; // @[MyOperators.scala 13:14:@16.4]
endmodule
