module Max3( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  input  [15:0] io_in1, // @[:@6.4]
  input  [15:0] io_in2, // @[:@6.4]
  input  [15:0] io_in3, // @[:@6.4]
  output [15:0] io_out // @[:@6.4]
);
  wire  _T_13; // @[Max3.scala 12:15:@8.4]
  wire  _T_14; // @[Max3.scala 12:34:@9.4]
  wire  _T_15; // @[Max3.scala 12:24:@10.4]
  wire  _T_16; // @[Max3.scala 14:21:@15.6]
  wire  _T_17; // @[Max3.scala 14:40:@16.6]
  wire  _T_18; // @[Max3.scala 14:30:@17.6]
  wire [15:0] _GEN_0; // @[Max3.scala 14:50:@18.6]
  assign _T_13 = io_in1 > io_in2; // @[Max3.scala 12:15:@8.4]
  assign _T_14 = io_in1 > io_in3; // @[Max3.scala 12:34:@9.4]
  assign _T_15 = _T_13 & _T_14; // @[Max3.scala 12:24:@10.4]
  assign _T_16 = io_in2 > io_in1; // @[Max3.scala 14:21:@15.6]
  assign _T_17 = io_in2 > io_in3; // @[Max3.scala 14:40:@16.6]
  assign _T_18 = _T_16 & _T_17; // @[Max3.scala 14:30:@17.6]
  assign _GEN_0 = _T_18 ? io_in2 : io_in3; // @[Max3.scala 14:50:@18.6]
  assign io_out = _T_15 ? io_in1 : _GEN_0; // @[Max3.scala 13:12:@12.6 Max3.scala 15:12:@19.8 Max3.scala 17:12:@22.8]
endmodule
