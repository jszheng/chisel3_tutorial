module VecShiftRegisterParam( // @[:@3.2]
  input        clock, // @[:@4.4]
  input        reset, // @[:@5.4]
  input  [7:0] io_in, // @[:@6.4]
  output [7:0] io_out // @[:@6.4]
);
  reg [7:0] delays_0; // @[VecShiftRegisterParam.scala 16:23:@19.4]
  reg [31:0] _RAND_0;
  reg [7:0] delays_1; // @[VecShiftRegisterParam.scala 16:23:@19.4]
  reg [31:0] _RAND_1;
  reg [7:0] delays_2; // @[VecShiftRegisterParam.scala 16:23:@19.4]
  reg [31:0] _RAND_2;
  reg [7:0] delays_3; // @[VecShiftRegisterParam.scala 16:23:@19.4]
  reg [31:0] _RAND_3;
  reg [7:0] delays_4; // @[VecShiftRegisterParam.scala 16:23:@19.4]
  reg [31:0] _RAND_4;
  reg [7:0] delays_5; // @[VecShiftRegisterParam.scala 16:23:@19.4]
  reg [31:0] _RAND_5;
  reg [7:0] delays_6; // @[VecShiftRegisterParam.scala 16:23:@19.4]
  reg [31:0] _RAND_6;
  reg [7:0] delays_7; // @[VecShiftRegisterParam.scala 16:23:@19.4]
  reg [31:0] _RAND_7;
  reg [7:0] delays_8; // @[VecShiftRegisterParam.scala 16:23:@19.4]
  reg [31:0] _RAND_8;
  reg [7:0] delays_9; // @[VecShiftRegisterParam.scala 16:23:@19.4]
  reg [31:0] _RAND_9;
  assign io_out = delays_9; // @[VecShiftRegisterParam.scala 23:10:@30.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  delays_0 = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  delays_1 = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  delays_2 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  delays_3 = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  delays_4 = _RAND_4[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  delays_5 = _RAND_5[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  delays_6 = _RAND_6[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  delays_7 = _RAND_7[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  delays_8 = _RAND_8[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  delays_9 = _RAND_9[7:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      delays_0 <= 8'h0;
    end else begin
      delays_0 <= io_in;
    end
    if (reset) begin
      delays_1 <= 8'h0;
    end else begin
      delays_1 <= delays_0;
    end
    if (reset) begin
      delays_2 <= 8'h0;
    end else begin
      delays_2 <= delays_1;
    end
    if (reset) begin
      delays_3 <= 8'h0;
    end else begin
      delays_3 <= delays_2;
    end
    if (reset) begin
      delays_4 <= 8'h0;
    end else begin
      delays_4 <= delays_3;
    end
    if (reset) begin
      delays_5 <= 8'h0;
    end else begin
      delays_5 <= delays_4;
    end
    if (reset) begin
      delays_6 <= 8'h0;
    end else begin
      delays_6 <= delays_5;
    end
    if (reset) begin
      delays_7 <= 8'h0;
    end else begin
      delays_7 <= delays_6;
    end
    if (reset) begin
      delays_8 <= 8'h0;
    end else begin
      delays_8 <= delays_7;
    end
    if (reset) begin
      delays_9 <= 8'h0;
    end else begin
      delays_9 <= delays_8;
    end
  end
endmodule
